
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER
-- DATE: Thu May 24 09:52:20 2018

	signal mem : ram_t := (
	

--			***** COLOR PALLETE *****


		0 =>	x"00000000", -- R: 0 G: 0 B: 0
		1 =>	x"00277FFF", -- R: 255 G: 127 B: 39
		2 =>	x"00383048", -- R: 72 G: 48 B: 56
		3 =>	x"0000E8B6", -- R: 182 G: 232 B: 0
		4 =>	x"00470000", -- R: 0 G: 0 B: 71
		5 =>	x"00700073", -- R: 115 G: 0 B: 112
		6 =>	x"00002D00", -- R: 0 G: 45 B: 0
		7 =>	x"0070006C", -- R: 108 G: 0 B: 112
		8 =>	x"00006F00", -- R: 0 G: 111 B: 0
		9 =>	x"00630000", -- R: 0 G: 0 B: 99
		10 =>	x"00007100", -- R: 0 G: 113 B: 0
		11 =>	x"0063006D", -- R: 109 G: 0 B: 99
		12 =>	x"000030BA", -- R: 186 G: 48 B: 0
		13 =>	x"00353B46", -- R: 70 G: 59 B: 53
		14 =>	x"007A0000", -- R: 0 G: 0 B: 122
		15 =>	x"006C002D", -- R: 45 G: 0 B: 108
		16 =>	x"00005300", -- R: 0 G: 83 B: 0
		17 =>	x"00490000", -- R: 0 G: 0 B: 73
		18 =>	x"00007400", -- R: 0 G: 116 B: 0
		19 =>	x"0068002D", -- R: 45 G: 0 B: 104
		20 =>	x"00005400", -- R: 0 G: 84 B: 0
		21 =>	x"00480000", -- R: 0 G: 0 B: 72
		22 =>	x"00007500", -- R: 0 G: 117 B: 0
		23 =>	x"006B002D", -- R: 45 G: 0 B: 107
		24 =>	x"00005500", -- R: 0 G: 85 B: 0
		25 =>	x"00410000", -- R: 0 G: 0 B: 65
		26 =>	x"00006600", -- R: 0 G: 102 B: 0
		27 =>	x"0079002D", -- R: 45 G: 0 B: 121
		28 =>	x"00004E00", -- R: 0 G: 78 B: 0
		29 =>	x"004C0000", -- R: 0 G: 0 B: 76
		30 =>	x"0072006F", -- R: 111 G: 0 B: 114
		31 =>	x"0052004F", -- R: 79 G: 0 B: 82
		32 =>	x"00730072", -- R: 114 G: 0 B: 115
		33 =>	x"004C0061", -- R: 97 G: 0 B: 76
		34 =>	x"006E002D", -- R: 45 G: 0 B: 110
		35 =>	x"00004300", -- R: 0 G: 67 B: 0
		36 =>	x"00530000", -- R: 0 G: 0 B: 83
		37 =>	x"00007300", -- R: 0 G: 115 B: 0
		38 =>	x"004B0000", -- R: 0 G: 0 B: 75
		39 =>	x"00680072", -- R: 114 G: 0 B: 104
		40 =>	x"00480052", -- R: 82 G: 0 B: 72
		41 =>	x"00650074", -- R: 116 G: 0 B: 101
		42 =>	x"00450045", -- R: 69 G: 0 B: 69
		43 =>	x"006C0076", -- R: 118 G: 0 B: 108
		44 =>	x"004C0056", -- R: 86 G: 0 B: 76
		45 =>	x"006C0074", -- R: 116 G: 0 B: 108
		46 =>	x"004C0054", -- R: 84 G: 0 B: 76
		47 =>	x"00720075", -- R: 117 G: 0 B: 114
		48 =>	x"00520055", -- R: 85 G: 0 B: 82
		49 =>	x"00730076", -- R: 118 G: 0 B: 115
		50 =>	x"00530045", -- R: 69 G: 0 B: 83
		51 =>	x"00740072", -- R: 114 G: 0 B: 116
		52 =>	x"00540052", -- R: 82 G: 0 B: 84
		53 =>	x"00620067", -- R: 103 G: 0 B: 98
		54 =>	x"00420047", -- R: 71 G: 0 B: 66
		55 =>	x"006E006C", -- R: 108 G: 0 B: 110
		56 =>	x"004E004C", -- R: 76 G: 0 B: 78
		57 =>	x"006E0062", -- R: 98 G: 0 B: 110
		58 =>	x"004E004F", -- R: 79 G: 0 B: 78
		59 =>	x"0050004C", -- R: 76 G: 0 B: 80
		60 =>	x"00700074", -- R: 116 G: 0 B: 112
		61 =>	x"00500054", -- R: 84 G: 0 B: 80
		62 =>	x"00680075", -- R: 117 G: 0 B: 104
		63 =>	x"00480055", -- R: 85 G: 0 B: 72
		64 =>	x"00690074", -- R: 116 G: 0 B: 105
		65 =>	x"00490054", -- R: 84 G: 0 B: 73
		66 =>	x"006A0061", -- R: 97 G: 0 B: 106
		67 =>	x"004A0050", -- R: 80 G: 0 B: 74
		68 =>	x"006B006F", -- R: 111 G: 0 B: 107
		69 =>	x"004B0052", -- R: 82 G: 0 B: 75
		70 =>	x"00660069", -- R: 105 G: 0 B: 102
		71 =>	x"00460049", -- R: 73 G: 0 B: 70
		72 =>	x"00660072", -- R: 114 G: 0 B: 102
		73 =>	x"00460052", -- R: 82 G: 0 B: 70
		74 =>	x"00640065", -- R: 101 G: 0 B: 100
		75 =>	x"00440045", -- R: 69 G: 0 B: 68
		76 =>	x"00680065", -- R: 101 G: 0 B: 104
		77 =>	x"0049004C", -- R: 76 G: 0 B: 73
		78 =>	x"00630073", -- R: 115 G: 0 B: 99
		79 =>	x"0043005A", -- R: 90 G: 0 B: 67
		80 =>	x"00640061", -- R: 97 G: 0 B: 100
		81 =>	x"0044004B", -- R: 75 G: 0 B: 68
		82 =>	x"0065006C", -- R: 108 G: 0 B: 101
		83 =>	x"00470052", -- R: 82 G: 0 B: 71
		84 =>	x"00650073", -- R: 115 G: 0 B: 101
		85 =>	x"00450053", -- R: 83 G: 0 B: 69
		86 =>	x"00420052", -- R: 82 G: 0 B: 66
		87 =>	x"007A0068", -- R: 104 G: 0 B: 122
		88 =>	x"00540057", -- R: 87 G: 0 B: 84
		89 =>	x"0043004E", -- R: 78 G: 0 B: 67
		90 =>	x"0048004B", -- R: 75 G: 0 B: 72
		91 =>	x"0043004C", -- R: 76 G: 0 B: 67
		92 =>	x"000042BB", -- R: 187 G: 66 B: 0
		93 =>	x"00344974", -- R: 116 G: 73 B: 52
		94 =>	x"007A0008", -- R: 8 G: 0 B: 122
		95 =>	x"0065006E", -- R: 110 G: 0 B: 101
		96 =>	x"00550053", -- R: 83 G: 0 B: 85
		97 =>	x"00610072", -- R: 114 G: 0 B: 97
		98 =>	x"00530041", -- R: 65 G: 0 B: 83
		99 =>	x"00310036", -- R: 54 G: 0 B: 49
		100 =>	x"00005C00", -- R: 0 G: 92 B: 0
		101 =>	x"002A002E", -- R: 46 G: 0 B: 42
		102 =>	x"00006200", -- R: 0 G: 98 B: 0
		103 =>	x"006D0070", -- R: 112 G: 0 B: 109
		104 =>	x"004C003B", -- R: 59 G: 0 B: 76
		105 =>	x"00050000", -- R: 0 G: 0 B: 5
		106 =>	x"0005627A", -- R: 122 G: 98 B: 5
		107 =>	x"000000E8", -- R: 232 G: 0 B: 0
		108 =>	x"00B64700", -- R: 0 G: 71 B: 182
		109 =>	x"00C40043", -- R: 67 G: 0 B: 196
		110 =>	x"00FDFDFD", -- R: 253 G: 253 B: 253
		111 =>	x"00FD6500", -- R: 0 G: 101 B: 253
		112 =>	x"005F0070", -- R: 112 G: 0 B: 95
		113 =>	x"00BB357A", -- R: 122 G: 53 B: 187
		114 =>	x"007F7A00", -- R: 0 G: 122 B: 127
		115 =>	x"004700C4", -- R: 196 G: 0 B: 71
		116 =>	x"00680069", -- R: 105 G: 0 B: 104
		117 =>	x"00006300", -- R: 0 G: 99 B: 0
		118 =>	x"00530074", -- R: 116 G: 0 B: 83
		119 =>	x"00660066", -- R: 102 G: 0 B: 102
		120 =>	x"00007800", -- R: 0 G: 120 B: 0
		121 =>	x"004798FF", -- R: 255 G: 152 B: 71
		122 =>	x"00FF0000", -- R: 0 G: 0 B: 255
		123 =>	x"0000FFFF", -- R: 255 G: 255 B: 0
		124 =>	x"000000FF", -- R: 255 G: 0 B: 0
		125 =>	x"00007F00", -- R: 0 G: 127 B: 0
		126 =>	x"004C4C4C", -- R: 76 G: 76 B: 76
		127 =>	x"007F007F", -- R: 127 G: 0 B: 127
		128 =>	x"0000007F", -- R: 127 G: 0 B: 0
		129 =>	x"00007F82", -- R: 130 G: 127 B: 0
		130 =>	x"00666666", -- R: 102 G: 102 B: 102
		131 =>	x"009800FF", -- R: 255 G: 0 B: 152
		132 =>	x"009800A4", -- R: 164 G: 0 B: 152
		133 =>	x"00980000", -- R: 0 G: 0 B: 152
		134 =>	x"005480D7", -- R: 215 G: 128 B: 84
		135 =>	x"00862138", -- R: 56 G: 33 B: 134
		136 =>	x"00990000", -- R: 0 G: 0 B: 153
		137 =>	x"00862136", -- R: 54 G: 33 B: 134
		138 =>	x"00980124", -- R: 36 G: 1 B: 152
		139 =>	x"00980095", -- R: 149 G: 0 B: 152
		140 =>	x"009800A5", -- R: 165 G: 0 B: 152
		141 =>	x"00980094", -- R: 148 G: 0 B: 152
		142 =>	x"009800DF", -- R: 223 G: 0 B: 152
		143 =>	x"009800A7", -- R: 167 G: 0 B: 152
		144 =>	x"0098016B", -- R: 107 G: 1 B: 152
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused
		255 =>	x"00000000", -- Unused

--			***** 16x16 IMAGES *****


		256 =>	x"01010101", -- IMG_16x16_background
		257 =>	x"01010101",
		258 =>	x"01010101",
		259 =>	x"01010101",
		260 =>	x"01010101",
		261 =>	x"01010101",
		262 =>	x"01010101",
		263 =>	x"01010101",
		264 =>	x"01010101",
		265 =>	x"01010101",
		266 =>	x"01010101",
		267 =>	x"01010101",
		268 =>	x"01010101",
		269 =>	x"01010101",
		270 =>	x"01010101",
		271 =>	x"01010101",
		272 =>	x"01010101",
		273 =>	x"01010101",
		274 =>	x"01010101",
		275 =>	x"01010101",
		276 =>	x"01010101",
		277 =>	x"01010101",
		278 =>	x"01010101",
		279 =>	x"01010101",
		280 =>	x"01010101",
		281 =>	x"01010101",
		282 =>	x"01010101",
		283 =>	x"01010101",
		284 =>	x"01010101",
		285 =>	x"01010101",
		286 =>	x"01010101",
		287 =>	x"01010101",
		288 =>	x"01010101",
		289 =>	x"01010101",
		290 =>	x"01010101",
		291 =>	x"01010101",
		292 =>	x"01010101",
		293 =>	x"01010101",
		294 =>	x"01010101",
		295 =>	x"01010101",
		296 =>	x"01010101",
		297 =>	x"01010101",
		298 =>	x"01010101",
		299 =>	x"01010101",
		300 =>	x"01010101",
		301 =>	x"01010101",
		302 =>	x"01010101",
		303 =>	x"01010101",
		304 =>	x"01010101",
		305 =>	x"01010101",
		306 =>	x"01010101",
		307 =>	x"01010101",
		308 =>	x"01010101",
		309 =>	x"01010101",
		310 =>	x"01010101",
		311 =>	x"01010101",
		312 =>	x"01010101",
		313 =>	x"01010101",
		314 =>	x"01010101",
		315 =>	x"01010101",
		316 =>	x"01010101",
		317 =>	x"01010101",
		318 =>	x"01010101",
		319 =>	x"01010101",
		320 =>	x"00000000", -- IMG_16x16_bang
		321 =>	x"00000000",
		322 =>	x"00000000",
		323 =>	x"00000000",
		324 =>	x"00000000",
		325 =>	x"00000000",
		326 =>	x"00000000",
		327 =>	x"00000000",
		328 =>	x"02030400",
		329 =>	x"00000000",
		330 =>	x"00000000",
		331 =>	x"00000000",
		332 =>	x"05060708",
		333 =>	x"090A0506",
		334 =>	x"07080B00",
		335 =>	x"000C0D0E",
		336 =>	x"0F101112",
		337 =>	x"13141516",
		338 =>	x"1718191A",
		339 =>	x"1B1C1D0A",
		340 =>	x"1E061F00",
		341 =>	x"20062112",
		342 =>	x"22232425",
		343 =>	x"17102625",
		344 =>	x"27062800",
		345 =>	x"29062A00",
		346 =>	x"2B062C00",
		347 =>	x"2D062E00",
		348 =>	x"2F063000",
		349 =>	x"31063200",
		350 =>	x"33063400",
		351 =>	x"35063600",
		352 =>	x"37063800",
		353 =>	x"39063A00",
		354 =>	x"07063B00",
		355 =>	x"3C063D00",
		356 =>	x"3E063F00",
		357 =>	x"40064100",
		358 =>	x"42064300",
		359 =>	x"44064500",
		360 =>	x"46064700",
		361 =>	x"48064900",
		362 =>	x"4A064B00",
		363 =>	x"4C064D00",
		364 =>	x"4E064F00",
		365 =>	x"50065100",
		366 =>	x"52065300",
		367 =>	x"54065500",
		368 =>	x"3C065600",
		369 =>	x"57065800",
		370 =>	x"57065900",
		371 =>	x"57065A00",
		372 =>	x"07080B00",
		373 =>	x"5B5C5D5E",
		374 =>	x"5F066000",
		375 =>	x"61066200",
		376 =>	x"63646566",
		377 =>	x"6700680A",
		378 =>	x"696A6B6C",
		379 =>	x"6D0A0506",
		380 =>	x"6E6F7071",
		381 =>	x"72037323",
		382 =>	x"74757616",
		383 =>	x"77646378",
		384 =>	x"79797979", -- IMG_16x16_car_blue
		385 =>	x"79797979",
		386 =>	x"79797979",
		387 =>	x"79797979",
		388 =>	x"79790000",
		389 =>	x"00797979",
		390 =>	x"79797979",
		391 =>	x"79797979",
		392 =>	x"79790000",
		393 =>	x"0079797A",
		394 =>	x"79797979",
		395 =>	x"79797979",
		396 =>	x"79797900",
		397 =>	x"7979797A",
		398 =>	x"7A797979",
		399 =>	x"79797979",
		400 =>	x"79797A7A",
		401 =>	x"7A7A7A7A",
		402 =>	x"7A7A7979",
		403 =>	x"00000079",
		404 =>	x"7900007A",
		405 =>	x"7A7A7A7A",
		406 =>	x"7A7A7A7A",
		407 =>	x"00000079",
		408 =>	x"79000000",
		409 =>	x"007B7B7B",
		410 =>	x"7A7A7A7A",
		411 =>	x"79007979",
		412 =>	x"79797A7A",
		413 =>	x"7A7B7B7B",
		414 =>	x"7B7A7A7A",
		415 =>	x"7A7A7A79",
		416 =>	x"79797A7A",
		417 =>	x"7A7B7B7B",
		418 =>	x"7B7A7A7A",
		419 =>	x"7A7A7A79",
		420 =>	x"79000000",
		421 =>	x"007B7B7B",
		422 =>	x"7A7A7A7A",
		423 =>	x"79007979",
		424 =>	x"7900007A",
		425 =>	x"7A7A7A7A",
		426 =>	x"7A7A7A7A",
		427 =>	x"00000079",
		428 =>	x"79797A7A",
		429 =>	x"7A7A7A7A",
		430 =>	x"7A7A7979",
		431 =>	x"00000079",
		432 =>	x"79797900",
		433 =>	x"7979797A",
		434 =>	x"7A797979",
		435 =>	x"79797979",
		436 =>	x"79790000",
		437 =>	x"0079797A",
		438 =>	x"79797979",
		439 =>	x"79797979",
		440 =>	x"79790000",
		441 =>	x"00797979",
		442 =>	x"79797979",
		443 =>	x"79797979",
		444 =>	x"79797979",
		445 =>	x"79797979",
		446 =>	x"79797979",
		447 =>	x"79797979",
		448 =>	x"79797979", -- IMG_16x16_car_red
		449 =>	x"79797979",
		450 =>	x"79797979",
		451 =>	x"79797979",
		452 =>	x"79790000",
		453 =>	x"00797979",
		454 =>	x"79797979",
		455 =>	x"79797979",
		456 =>	x"79790000",
		457 =>	x"0079797C",
		458 =>	x"79797979",
		459 =>	x"79797979",
		460 =>	x"79797900",
		461 =>	x"7979797C",
		462 =>	x"7C797979",
		463 =>	x"79797979",
		464 =>	x"79797C7C",
		465 =>	x"7C7C7C7C",
		466 =>	x"7C7C7979",
		467 =>	x"00000079",
		468 =>	x"7900007C",
		469 =>	x"7C7C7C7C",
		470 =>	x"7C7C7C7C",
		471 =>	x"00000079",
		472 =>	x"79000000",
		473 =>	x"007B7B7B",
		474 =>	x"7C7C7C7C",
		475 =>	x"79007979",
		476 =>	x"79797C7C",
		477 =>	x"7C7B7B7B",
		478 =>	x"7B7C7C7C",
		479 =>	x"7C7C7C79",
		480 =>	x"79797C7C",
		481 =>	x"7C7B7B7B",
		482 =>	x"7B7C7C7C",
		483 =>	x"7C7C7C79",
		484 =>	x"79000000",
		485 =>	x"007B7B7B",
		486 =>	x"7C7C7C7C",
		487 =>	x"79007979",
		488 =>	x"7900007C",
		489 =>	x"7C7C7C7C",
		490 =>	x"7C7C7C7C",
		491 =>	x"00000079",
		492 =>	x"79797C7C",
		493 =>	x"7C7C7C7C",
		494 =>	x"7C7C7979",
		495 =>	x"00000079",
		496 =>	x"79797900",
		497 =>	x"7979797C",
		498 =>	x"7C797979",
		499 =>	x"79797979",
		500 =>	x"79790000",
		501 =>	x"0079797C",
		502 =>	x"79797979",
		503 =>	x"79797979",
		504 =>	x"79790000",
		505 =>	x"00797979",
		506 =>	x"79797979",
		507 =>	x"79797979",
		508 =>	x"79797979",
		509 =>	x"79797979",
		510 =>	x"79797979",
		511 =>	x"79797979",
		512 =>	x"01010101", -- IMG_16x16_flag
		513 =>	x"01010101",
		514 =>	x"01010101",
		515 =>	x"01010101",
		516 =>	x"01017B7B",
		517 =>	x"01010101",
		518 =>	x"01010101",
		519 =>	x"01010101",
		520 =>	x"01017B7B",
		521 =>	x"7B7B0101",
		522 =>	x"01010101",
		523 =>	x"01010101",
		524 =>	x"01017B7B",
		525 =>	x"7B7B7B7B",
		526 =>	x"01010101",
		527 =>	x"01010101",
		528 =>	x"01017B7B",
		529 =>	x"7B7B7B7B",
		530 =>	x"7B7B0101",
		531 =>	x"01010101",
		532 =>	x"01017B7B",
		533 =>	x"7B7B7B7B",
		534 =>	x"7B7B7B7B",
		535 =>	x"01010101",
		536 =>	x"01017B7B",
		537 =>	x"7B7B7B7B",
		538 =>	x"7B7B0101",
		539 =>	x"01010101",
		540 =>	x"01017B7B",
		541 =>	x"7B7B7B7B",
		542 =>	x"01010101",
		543 =>	x"01010101",
		544 =>	x"01017B7B",
		545 =>	x"7B7B0101",
		546 =>	x"01010101",
		547 =>	x"01010101",
		548 =>	x"01017B7B",
		549 =>	x"01010101",
		550 =>	x"01010101",
		551 =>	x"01010101",
		552 =>	x"01017B7B",
		553 =>	x"01010101",
		554 =>	x"01010101",
		555 =>	x"01010101",
		556 =>	x"01017B7B",
		557 =>	x"01010101",
		558 =>	x"01010101",
		559 =>	x"01010101",
		560 =>	x"01017B7B",
		561 =>	x"01010101",
		562 =>	x"01010101",
		563 =>	x"01010101",
		564 =>	x"017B7B7B",
		565 =>	x"7B010101",
		566 =>	x"01010101",
		567 =>	x"01010101",
		568 =>	x"017B7B7B",
		569 =>	x"7B010101",
		570 =>	x"01010101",
		571 =>	x"01010101",
		572 =>	x"01010101",
		573 =>	x"01010101",
		574 =>	x"01010101",
		575 =>	x"01010101",
		576 =>	x"7D7D7D7D", -- IMG_16x16_map_element_00
		577 =>	x"7D7D7E7D",
		578 =>	x"7E7E7D7D",
		579 =>	x"7D7D7D7D",
		580 =>	x"7D7D7D7D",
		581 =>	x"7F80807F",
		582 =>	x"807F807E",
		583 =>	x"7D7D7D7D",
		584 =>	x"7D7D7E80",
		585 =>	x"7F80807F",
		586 =>	x"81828080",
		587 =>	x"7D7D7D7D",
		588 =>	x"7D7D7F80",
		589 =>	x"80807F7F",
		590 =>	x"80807F7F",
		591 =>	x"80807D7D",
		592 =>	x"7D7E8080",
		593 =>	x"80807F7F",
		594 =>	x"807C7F7F",
		595 =>	x"7F7E7E7D",
		596 =>	x"7E7F7F80",
		597 =>	x"807C7F7F",
		598 =>	x"807C7F80",
		599 =>	x"8080807E",
		600 =>	x"7E808080",
		601 =>	x"8080807F",
		602 =>	x"8080807C",
		603 =>	x"7C80807E",
		604 =>	x"7E817F7F",
		605 =>	x"807F7F7E",
		606 =>	x"7F7F807F",
		607 =>	x"7C807E7E",
		608 =>	x"7E808081",
		609 =>	x"80808080",
		610 =>	x"8080807C",
		611 =>	x"8080807E",
		612 =>	x"7E808080",
		613 =>	x"8081807F",
		614 =>	x"80807F80",
		615 =>	x"7F807F7E",
		616 =>	x"7E7F8080",
		617 =>	x"80807F80",
		618 =>	x"7C7F8080",
		619 =>	x"7F7E7F7E",
		620 =>	x"7D80807F",
		621 =>	x"7F7F7F80",
		622 =>	x"807F7F80",
		623 =>	x"7F7F7E7D",
		624 =>	x"7D7D7F80",
		625 =>	x"807F8080",
		626 =>	x"7F7F7F80",
		627 =>	x"80807E7D",
		628 =>	x"7D7D7E81",
		629 =>	x"807F8180",
		630 =>	x"7F7F8080",
		631 =>	x"7F7E7D7D",
		632 =>	x"7D7D7D7D",
		633 =>	x"7E808181",
		634 =>	x"807C7E7D",
		635 =>	x"7D7D7D7D",
		636 =>	x"7D7D7D7D",
		637 =>	x"7D7D7E7E",
		638 =>	x"7E7E7D7D",
		639 =>	x"7D7D7D7D",
		640 =>	x"83838383", -- IMG_16x16_map_element_01
		641 =>	x"83838383",
		642 =>	x"83838383",
		643 =>	x"83838485",
		644 =>	x"83838383",
		645 =>	x"83838383",
		646 =>	x"83838383",
		647 =>	x"83838485",
		648 =>	x"83838383",
		649 =>	x"83838383",
		650 =>	x"83838383",
		651 =>	x"83838485",
		652 =>	x"83838383",
		653 =>	x"83838383",
		654 =>	x"83838383",
		655 =>	x"83838485",
		656 =>	x"83838383",
		657 =>	x"83838383",
		658 =>	x"83838383",
		659 =>	x"83838485",
		660 =>	x"83838383",
		661 =>	x"83838383",
		662 =>	x"83838383",
		663 =>	x"83838485",
		664 =>	x"83838383",
		665 =>	x"83838383",
		666 =>	x"83838383",
		667 =>	x"83838485",
		668 =>	x"83838383",
		669 =>	x"83838383",
		670 =>	x"83838383",
		671 =>	x"83838485",
		672 =>	x"83838383",
		673 =>	x"83838383",
		674 =>	x"83838383",
		675 =>	x"83838485",
		676 =>	x"83838383",
		677 =>	x"83838383",
		678 =>	x"83838383",
		679 =>	x"83838485",
		680 =>	x"83838383",
		681 =>	x"83838383",
		682 =>	x"83838383",
		683 =>	x"83838485",
		684 =>	x"83838383",
		685 =>	x"83838383",
		686 =>	x"83838383",
		687 =>	x"83838485",
		688 =>	x"83838383",
		689 =>	x"83838383",
		690 =>	x"83838383",
		691 =>	x"83838485",
		692 =>	x"83838383",
		693 =>	x"83838383",
		694 =>	x"83838383",
		695 =>	x"83838485",
		696 =>	x"83838383",
		697 =>	x"83838383",
		698 =>	x"83838383",
		699 =>	x"83838485",
		700 =>	x"83838383",
		701 =>	x"83838383",
		702 =>	x"83838383",
		703 =>	x"83838485",
		704 =>	x"86878885", -- IMG_16x16_map_element_02
		705 =>	x"85858585",
		706 =>	x"85858585",
		707 =>	x"85858585",
		708 =>	x"898A8B8C",
		709 =>	x"84848484",
		710 =>	x"84848484",
		711 =>	x"84848484",
		712 =>	x"888D8383",
		713 =>	x"83838383",
		714 =>	x"83838383",
		715 =>	x"83838383",
		716 =>	x"85848383",
		717 =>	x"83838383",
		718 =>	x"83838383",
		719 =>	x"83838383",
		720 =>	x"85848383",
		721 =>	x"83838383",
		722 =>	x"83838383",
		723 =>	x"83838383",
		724 =>	x"85848383",
		725 =>	x"83838383",
		726 =>	x"83838383",
		727 =>	x"83838383",
		728 =>	x"85848383",
		729 =>	x"83838383",
		730 =>	x"83838383",
		731 =>	x"83838383",
		732 =>	x"85848383",
		733 =>	x"83838383",
		734 =>	x"83838383",
		735 =>	x"83838383",
		736 =>	x"85848383",
		737 =>	x"83838383",
		738 =>	x"83838383",
		739 =>	x"83838383",
		740 =>	x"85848383",
		741 =>	x"83838383",
		742 =>	x"83838383",
		743 =>	x"83838383",
		744 =>	x"85848383",
		745 =>	x"83838383",
		746 =>	x"83838383",
		747 =>	x"83838383",
		748 =>	x"85848383",
		749 =>	x"83838383",
		750 =>	x"83838383",
		751 =>	x"83838383",
		752 =>	x"85848383",
		753 =>	x"83838383",
		754 =>	x"83838383",
		755 =>	x"83838383",
		756 =>	x"888D8383",
		757 =>	x"83838383",
		758 =>	x"83838383",
		759 =>	x"83838383",
		760 =>	x"898A8B8C",
		761 =>	x"84848484",
		762 =>	x"84848484",
		763 =>	x"84848484",
		764 =>	x"86878885",
		765 =>	x"85858585",
		766 =>	x"85858585",
		767 =>	x"85858585",
		768 =>	x"85848383", -- IMG_16x16_map_element_03
		769 =>	x"83838383",
		770 =>	x"83838383",
		771 =>	x"83838485",
		772 =>	x"848E8383",
		773 =>	x"83838383",
		774 =>	x"83838383",
		775 =>	x"83838E84",
		776 =>	x"83838383",
		777 =>	x"83838383",
		778 =>	x"83838383",
		779 =>	x"83838383",
		780 =>	x"83838383",
		781 =>	x"83838383",
		782 =>	x"83838383",
		783 =>	x"83838383",
		784 =>	x"83838383",
		785 =>	x"83838383",
		786 =>	x"83838383",
		787 =>	x"83838383",
		788 =>	x"83838383",
		789 =>	x"83838383",
		790 =>	x"83838383",
		791 =>	x"83838383",
		792 =>	x"83838383",
		793 =>	x"83838383",
		794 =>	x"83838383",
		795 =>	x"83838383",
		796 =>	x"83838383",
		797 =>	x"83838383",
		798 =>	x"83838383",
		799 =>	x"83838383",
		800 =>	x"83838383",
		801 =>	x"83838383",
		802 =>	x"83838383",
		803 =>	x"83838383",
		804 =>	x"83838383",
		805 =>	x"83838383",
		806 =>	x"83838383",
		807 =>	x"83838383",
		808 =>	x"83838383",
		809 =>	x"83838383",
		810 =>	x"83838383",
		811 =>	x"83838383",
		812 =>	x"83838383",
		813 =>	x"83838383",
		814 =>	x"83838383",
		815 =>	x"83838383",
		816 =>	x"83838383",
		817 =>	x"83838383",
		818 =>	x"83838383",
		819 =>	x"83838383",
		820 =>	x"83838383",
		821 =>	x"83838383",
		822 =>	x"83838383",
		823 =>	x"83838383",
		824 =>	x"848E8383",
		825 =>	x"83838383",
		826 =>	x"83838383",
		827 =>	x"83838E84",
		828 =>	x"85848383",
		829 =>	x"83838383",
		830 =>	x"83838383",
		831 =>	x"83838485",
		832 =>	x"85858585", -- IMG_16x16_map_element_04
		833 =>	x"85858585",
		834 =>	x"85858585",
		835 =>	x"85888786",
		836 =>	x"84848484",
		837 =>	x"84848484",
		838 =>	x"84848484",
		839 =>	x"8C8B8A89",
		840 =>	x"83838383",
		841 =>	x"83838383",
		842 =>	x"83838383",
		843 =>	x"83838D88",
		844 =>	x"83838383",
		845 =>	x"83838383",
		846 =>	x"83838383",
		847 =>	x"83838485",
		848 =>	x"83838383",
		849 =>	x"83838383",
		850 =>	x"83838383",
		851 =>	x"83838485",
		852 =>	x"83838383",
		853 =>	x"83838383",
		854 =>	x"83838383",
		855 =>	x"83838485",
		856 =>	x"83838383",
		857 =>	x"83838383",
		858 =>	x"83838383",
		859 =>	x"83838485",
		860 =>	x"83838383",
		861 =>	x"83838383",
		862 =>	x"83838383",
		863 =>	x"83838485",
		864 =>	x"83838383",
		865 =>	x"83838383",
		866 =>	x"83838383",
		867 =>	x"83838485",
		868 =>	x"83838383",
		869 =>	x"83838383",
		870 =>	x"83838383",
		871 =>	x"83838485",
		872 =>	x"83838383",
		873 =>	x"83838383",
		874 =>	x"83838383",
		875 =>	x"83838485",
		876 =>	x"83838383",
		877 =>	x"83838383",
		878 =>	x"83838383",
		879 =>	x"83838485",
		880 =>	x"83838383",
		881 =>	x"83838383",
		882 =>	x"83838383",
		883 =>	x"83838485",
		884 =>	x"83838383",
		885 =>	x"83838383",
		886 =>	x"83838383",
		887 =>	x"83838D88",
		888 =>	x"84848484",
		889 =>	x"84848484",
		890 =>	x"84848484",
		891 =>	x"8C8B8A89",
		892 =>	x"85858585",
		893 =>	x"85858585",
		894 =>	x"85858585",
		895 =>	x"85888786",
		896 =>	x"85848383", -- IMG_16x16_map_element_05
		897 =>	x"83838383",
		898 =>	x"83838383",
		899 =>	x"83838383",
		900 =>	x"85848383",
		901 =>	x"83838383",
		902 =>	x"83838383",
		903 =>	x"83838383",
		904 =>	x"85848383",
		905 =>	x"83838383",
		906 =>	x"83838383",
		907 =>	x"83838383",
		908 =>	x"85848383",
		909 =>	x"83838383",
		910 =>	x"83838383",
		911 =>	x"83838383",
		912 =>	x"85848383",
		913 =>	x"83838383",
		914 =>	x"83838383",
		915 =>	x"83838383",
		916 =>	x"85848383",
		917 =>	x"83838383",
		918 =>	x"83838383",
		919 =>	x"83838383",
		920 =>	x"85848383",
		921 =>	x"83838383",
		922 =>	x"83838383",
		923 =>	x"83838383",
		924 =>	x"85848383",
		925 =>	x"83838383",
		926 =>	x"83838383",
		927 =>	x"83838383",
		928 =>	x"85848383",
		929 =>	x"83838383",
		930 =>	x"83838383",
		931 =>	x"83838383",
		932 =>	x"85848383",
		933 =>	x"83838383",
		934 =>	x"83838383",
		935 =>	x"83838383",
		936 =>	x"85848383",
		937 =>	x"83838383",
		938 =>	x"83838383",
		939 =>	x"83838383",
		940 =>	x"85848383",
		941 =>	x"83838383",
		942 =>	x"83838383",
		943 =>	x"83838383",
		944 =>	x"85848383",
		945 =>	x"83838383",
		946 =>	x"83838383",
		947 =>	x"83838383",
		948 =>	x"888D8383",
		949 =>	x"83838383",
		950 =>	x"83838383",
		951 =>	x"83838383",
		952 =>	x"898A8B8C",
		953 =>	x"84848484",
		954 =>	x"84848484",
		955 =>	x"84848484",
		956 =>	x"86878885",
		957 =>	x"85858585",
		958 =>	x"85858585",
		959 =>	x"85858585",
		960 =>	x"83838383", -- IMG_16x16_map_element_06
		961 =>	x"83838383",
		962 =>	x"83838383",
		963 =>	x"83838383",
		964 =>	x"83838383",
		965 =>	x"83838383",
		966 =>	x"83838383",
		967 =>	x"83838383",
		968 =>	x"83838383",
		969 =>	x"83838383",
		970 =>	x"83838383",
		971 =>	x"83838383",
		972 =>	x"83838383",
		973 =>	x"83838383",
		974 =>	x"83838383",
		975 =>	x"83838383",
		976 =>	x"83838383",
		977 =>	x"83838383",
		978 =>	x"83838383",
		979 =>	x"83838383",
		980 =>	x"83838383",
		981 =>	x"83838383",
		982 =>	x"83838383",
		983 =>	x"83838383",
		984 =>	x"83838383",
		985 =>	x"83838383",
		986 =>	x"83838383",
		987 =>	x"83838383",
		988 =>	x"83838383",
		989 =>	x"83838383",
		990 =>	x"83838383",
		991 =>	x"83838383",
		992 =>	x"83838383",
		993 =>	x"83838383",
		994 =>	x"83838383",
		995 =>	x"83838383",
		996 =>	x"83838383",
		997 =>	x"83838383",
		998 =>	x"83838383",
		999 =>	x"83838383",
		1000 =>	x"83838383",
		1001 =>	x"83838383",
		1002 =>	x"83838383",
		1003 =>	x"83838383",
		1004 =>	x"83838383",
		1005 =>	x"83838383",
		1006 =>	x"83838383",
		1007 =>	x"83838383",
		1008 =>	x"83838383",
		1009 =>	x"83838383",
		1010 =>	x"83838383",
		1011 =>	x"83838383",
		1012 =>	x"83838383",
		1013 =>	x"83838383",
		1014 =>	x"83838383",
		1015 =>	x"83838383",
		1016 =>	x"84848484",
		1017 =>	x"84848484",
		1018 =>	x"84848484",
		1019 =>	x"84848484",
		1020 =>	x"85858585",
		1021 =>	x"85858585",
		1022 =>	x"85858585",
		1023 =>	x"85858585",
		1024 =>	x"83838383", -- IMG_16x16_map_element_07
		1025 =>	x"83838383",
		1026 =>	x"83838383",
		1027 =>	x"83838485",
		1028 =>	x"83838383",
		1029 =>	x"83838383",
		1030 =>	x"83838383",
		1031 =>	x"83838485",
		1032 =>	x"83838383",
		1033 =>	x"83838383",
		1034 =>	x"83838383",
		1035 =>	x"83838485",
		1036 =>	x"83838383",
		1037 =>	x"83838383",
		1038 =>	x"83838383",
		1039 =>	x"83838485",
		1040 =>	x"83838383",
		1041 =>	x"83838383",
		1042 =>	x"83838383",
		1043 =>	x"83838485",
		1044 =>	x"83838383",
		1045 =>	x"83838383",
		1046 =>	x"83838383",
		1047 =>	x"83838485",
		1048 =>	x"83838383",
		1049 =>	x"83838383",
		1050 =>	x"83838383",
		1051 =>	x"83838485",
		1052 =>	x"83838383",
		1053 =>	x"83838383",
		1054 =>	x"83838383",
		1055 =>	x"83838485",
		1056 =>	x"83838383",
		1057 =>	x"83838383",
		1058 =>	x"83838383",
		1059 =>	x"83838485",
		1060 =>	x"83838383",
		1061 =>	x"83838383",
		1062 =>	x"83838383",
		1063 =>	x"83838485",
		1064 =>	x"83838383",
		1065 =>	x"83838383",
		1066 =>	x"83838383",
		1067 =>	x"83838485",
		1068 =>	x"83838383",
		1069 =>	x"83838383",
		1070 =>	x"83838383",
		1071 =>	x"83838485",
		1072 =>	x"83838383",
		1073 =>	x"83838383",
		1074 =>	x"83838383",
		1075 =>	x"83838485",
		1076 =>	x"83838383",
		1077 =>	x"83838383",
		1078 =>	x"83838383",
		1079 =>	x"83838D88",
		1080 =>	x"84848484",
		1081 =>	x"84848484",
		1082 =>	x"84848484",
		1083 =>	x"8C8B8A89",
		1084 =>	x"85858585",
		1085 =>	x"85858585",
		1086 =>	x"85858585",
		1087 =>	x"85888786",
		1088 =>	x"85848383", -- IMG_16x16_map_element_08
		1089 =>	x"83838383",
		1090 =>	x"83838383",
		1091 =>	x"83838485",
		1092 =>	x"85848383",
		1093 =>	x"83838383",
		1094 =>	x"83838383",
		1095 =>	x"83838E84",
		1096 =>	x"85848383",
		1097 =>	x"83838383",
		1098 =>	x"83838383",
		1099 =>	x"83838383",
		1100 =>	x"85848383",
		1101 =>	x"83838383",
		1102 =>	x"83838383",
		1103 =>	x"83838383",
		1104 =>	x"85848383",
		1105 =>	x"83838383",
		1106 =>	x"83838383",
		1107 =>	x"83838383",
		1108 =>	x"85848383",
		1109 =>	x"83838383",
		1110 =>	x"83838383",
		1111 =>	x"83838383",
		1112 =>	x"85848383",
		1113 =>	x"83838383",
		1114 =>	x"83838383",
		1115 =>	x"83838383",
		1116 =>	x"85848383",
		1117 =>	x"83838383",
		1118 =>	x"83838383",
		1119 =>	x"83838383",
		1120 =>	x"85848383",
		1121 =>	x"83838383",
		1122 =>	x"83838383",
		1123 =>	x"83838383",
		1124 =>	x"85848383",
		1125 =>	x"83838383",
		1126 =>	x"83838383",
		1127 =>	x"83838383",
		1128 =>	x"85848383",
		1129 =>	x"83838383",
		1130 =>	x"83838383",
		1131 =>	x"83838383",
		1132 =>	x"85848383",
		1133 =>	x"83838383",
		1134 =>	x"83838383",
		1135 =>	x"83838383",
		1136 =>	x"85848383",
		1137 =>	x"83838383",
		1138 =>	x"83838383",
		1139 =>	x"83838383",
		1140 =>	x"888D8383",
		1141 =>	x"83838383",
		1142 =>	x"83838383",
		1143 =>	x"83838383",
		1144 =>	x"898A8B8C",
		1145 =>	x"84848484",
		1146 =>	x"84848484",
		1147 =>	x"84848484",
		1148 =>	x"86878885",
		1149 =>	x"85858585",
		1150 =>	x"85858585",
		1151 =>	x"85858585",
		1152 =>	x"85848383", -- IMG_16x16_map_element_09
		1153 =>	x"83838383",
		1154 =>	x"83838383",
		1155 =>	x"83838485",
		1156 =>	x"85848383",
		1157 =>	x"83838383",
		1158 =>	x"83838383",
		1159 =>	x"83838485",
		1160 =>	x"85848383",
		1161 =>	x"83838383",
		1162 =>	x"83838383",
		1163 =>	x"83838485",
		1164 =>	x"85848383",
		1165 =>	x"83838383",
		1166 =>	x"83838383",
		1167 =>	x"83838485",
		1168 =>	x"85848383",
		1169 =>	x"83838383",
		1170 =>	x"83838383",
		1171 =>	x"83838485",
		1172 =>	x"85848383",
		1173 =>	x"83838383",
		1174 =>	x"83838383",
		1175 =>	x"83838485",
		1176 =>	x"85848383",
		1177 =>	x"83838383",
		1178 =>	x"83838383",
		1179 =>	x"83838485",
		1180 =>	x"85848383",
		1181 =>	x"83838383",
		1182 =>	x"83838383",
		1183 =>	x"83838485",
		1184 =>	x"85848383",
		1185 =>	x"83838383",
		1186 =>	x"83838383",
		1187 =>	x"83838485",
		1188 =>	x"85848383",
		1189 =>	x"83838383",
		1190 =>	x"83838383",
		1191 =>	x"83838485",
		1192 =>	x"85848383",
		1193 =>	x"83838383",
		1194 =>	x"83838383",
		1195 =>	x"83838485",
		1196 =>	x"85848383",
		1197 =>	x"83838383",
		1198 =>	x"83838383",
		1199 =>	x"83838485",
		1200 =>	x"85848383",
		1201 =>	x"83838383",
		1202 =>	x"83838383",
		1203 =>	x"83838485",
		1204 =>	x"888D8383",
		1205 =>	x"83838383",
		1206 =>	x"83838383",
		1207 =>	x"83838D88",
		1208 =>	x"898A8B8C",
		1209 =>	x"84848484",
		1210 =>	x"84848484",
		1211 =>	x"8C8B8A89",
		1212 =>	x"86878885",
		1213 =>	x"85858585",
		1214 =>	x"85858585",
		1215 =>	x"85888786",
		1216 =>	x"85848383", -- IMG_16x16_map_element_10
		1217 =>	x"83838383",
		1218 =>	x"83838383",
		1219 =>	x"83838485",
		1220 =>	x"848E8383",
		1221 =>	x"83838383",
		1222 =>	x"83838383",
		1223 =>	x"83838485",
		1224 =>	x"83838383",
		1225 =>	x"83838383",
		1226 =>	x"83838383",
		1227 =>	x"83838485",
		1228 =>	x"83838383",
		1229 =>	x"83838383",
		1230 =>	x"83838383",
		1231 =>	x"83838485",
		1232 =>	x"83838383",
		1233 =>	x"83838383",
		1234 =>	x"83838383",
		1235 =>	x"83838485",
		1236 =>	x"83838383",
		1237 =>	x"83838383",
		1238 =>	x"83838383",
		1239 =>	x"83838485",
		1240 =>	x"83838383",
		1241 =>	x"83838383",
		1242 =>	x"83838383",
		1243 =>	x"83838485",
		1244 =>	x"83838383",
		1245 =>	x"83838383",
		1246 =>	x"83838383",
		1247 =>	x"83838485",
		1248 =>	x"83838383",
		1249 =>	x"83838383",
		1250 =>	x"83838383",
		1251 =>	x"83838485",
		1252 =>	x"83838383",
		1253 =>	x"83838383",
		1254 =>	x"83838383",
		1255 =>	x"83838485",
		1256 =>	x"83838383",
		1257 =>	x"83838383",
		1258 =>	x"83838383",
		1259 =>	x"83838485",
		1260 =>	x"83838383",
		1261 =>	x"83838383",
		1262 =>	x"83838383",
		1263 =>	x"83838485",
		1264 =>	x"83838383",
		1265 =>	x"83838383",
		1266 =>	x"83838383",
		1267 =>	x"83838485",
		1268 =>	x"83838383",
		1269 =>	x"83838383",
		1270 =>	x"83838383",
		1271 =>	x"83838D88",
		1272 =>	x"84848484",
		1273 =>	x"84848484",
		1274 =>	x"84848484",
		1275 =>	x"8C8B8A89",
		1276 =>	x"85858585",
		1277 =>	x"85858585",
		1278 =>	x"85858585",
		1279 =>	x"85888786",
		1280 =>	x"86878885", -- IMG_16x16_map_element_11
		1281 =>	x"85858585",
		1282 =>	x"85858585",
		1283 =>	x"85858585",
		1284 =>	x"898A8B8C",
		1285 =>	x"84848484",
		1286 =>	x"84848484",
		1287 =>	x"84848484",
		1288 =>	x"888D8383",
		1289 =>	x"83838383",
		1290 =>	x"83838383",
		1291 =>	x"83838383",
		1292 =>	x"85848383",
		1293 =>	x"83838383",
		1294 =>	x"83838383",
		1295 =>	x"83838383",
		1296 =>	x"85848383",
		1297 =>	x"83838383",
		1298 =>	x"83838383",
		1299 =>	x"83838383",
		1300 =>	x"85848383",
		1301 =>	x"83838383",
		1302 =>	x"83838383",
		1303 =>	x"83838383",
		1304 =>	x"85848383",
		1305 =>	x"83838383",
		1306 =>	x"83838383",
		1307 =>	x"83838383",
		1308 =>	x"85848383",
		1309 =>	x"83838383",
		1310 =>	x"83838383",
		1311 =>	x"83838383",
		1312 =>	x"85848383",
		1313 =>	x"83838383",
		1314 =>	x"83838383",
		1315 =>	x"83838383",
		1316 =>	x"85848383",
		1317 =>	x"83838383",
		1318 =>	x"83838383",
		1319 =>	x"83838383",
		1320 =>	x"85848383",
		1321 =>	x"83838383",
		1322 =>	x"83838383",
		1323 =>	x"83838383",
		1324 =>	x"85848383",
		1325 =>	x"83838383",
		1326 =>	x"83838383",
		1327 =>	x"83838383",
		1328 =>	x"85848383",
		1329 =>	x"83838383",
		1330 =>	x"83838383",
		1331 =>	x"83838383",
		1332 =>	x"85848383",
		1333 =>	x"83838383",
		1334 =>	x"83838383",
		1335 =>	x"83838383",
		1336 =>	x"85848383",
		1337 =>	x"83838383",
		1338 =>	x"83838383",
		1339 =>	x"83838383",
		1340 =>	x"85848383",
		1341 =>	x"83838383",
		1342 =>	x"83838383",
		1343 =>	x"83838383",
		1344 =>	x"85858585", -- IMG_16x16_map_element_12
		1345 =>	x"85858585",
		1346 =>	x"85858585",
		1347 =>	x"85858585",
		1348 =>	x"84848484",
		1349 =>	x"84848484",
		1350 =>	x"84848484",
		1351 =>	x"84848484",
		1352 =>	x"83838383",
		1353 =>	x"83838383",
		1354 =>	x"83838383",
		1355 =>	x"83838383",
		1356 =>	x"83838383",
		1357 =>	x"83838383",
		1358 =>	x"83838383",
		1359 =>	x"83838383",
		1360 =>	x"83838383",
		1361 =>	x"83838383",
		1362 =>	x"83838383",
		1363 =>	x"83838383",
		1364 =>	x"83838383",
		1365 =>	x"83838383",
		1366 =>	x"83838383",
		1367 =>	x"83838383",
		1368 =>	x"83838383",
		1369 =>	x"83838383",
		1370 =>	x"83838383",
		1371 =>	x"83838383",
		1372 =>	x"83838383",
		1373 =>	x"83838383",
		1374 =>	x"83838383",
		1375 =>	x"83838383",
		1376 =>	x"83838383",
		1377 =>	x"83838383",
		1378 =>	x"83838383",
		1379 =>	x"83838383",
		1380 =>	x"83838383",
		1381 =>	x"83838383",
		1382 =>	x"83838383",
		1383 =>	x"83838383",
		1384 =>	x"83838383",
		1385 =>	x"83838383",
		1386 =>	x"83838383",
		1387 =>	x"83838383",
		1388 =>	x"83838383",
		1389 =>	x"83838383",
		1390 =>	x"83838383",
		1391 =>	x"83838383",
		1392 =>	x"83838383",
		1393 =>	x"83838383",
		1394 =>	x"83838383",
		1395 =>	x"83838383",
		1396 =>	x"83838383",
		1397 =>	x"83838383",
		1398 =>	x"83838383",
		1399 =>	x"83838383",
		1400 =>	x"848E8383",
		1401 =>	x"83838383",
		1402 =>	x"83838383",
		1403 =>	x"83838E84",
		1404 =>	x"85848383",
		1405 =>	x"83838383",
		1406 =>	x"83838383",
		1407 =>	x"83838485",
		1408 =>	x"85848383", -- IMG_16x16_map_element_13
		1409 =>	x"83838383",
		1410 =>	x"83838383",
		1411 =>	x"83838485",
		1412 =>	x"85848383",
		1413 =>	x"83838383",
		1414 =>	x"83838383",
		1415 =>	x"83838E84",
		1416 =>	x"85848383",
		1417 =>	x"83838383",
		1418 =>	x"83838383",
		1419 =>	x"83838383",
		1420 =>	x"85848383",
		1421 =>	x"83838383",
		1422 =>	x"83838383",
		1423 =>	x"83838383",
		1424 =>	x"85848383",
		1425 =>	x"83838383",
		1426 =>	x"83838383",
		1427 =>	x"83838383",
		1428 =>	x"85848383",
		1429 =>	x"83838383",
		1430 =>	x"83838383",
		1431 =>	x"83838383",
		1432 =>	x"85848383",
		1433 =>	x"83838383",
		1434 =>	x"83838383",
		1435 =>	x"83838383",
		1436 =>	x"85848383",
		1437 =>	x"83838383",
		1438 =>	x"83838383",
		1439 =>	x"83838383",
		1440 =>	x"85848383",
		1441 =>	x"83838383",
		1442 =>	x"83838383",
		1443 =>	x"83838383",
		1444 =>	x"85848383",
		1445 =>	x"83838383",
		1446 =>	x"83838383",
		1447 =>	x"83838383",
		1448 =>	x"85848383",
		1449 =>	x"83838383",
		1450 =>	x"83838383",
		1451 =>	x"83838383",
		1452 =>	x"85848383",
		1453 =>	x"83838383",
		1454 =>	x"83838383",
		1455 =>	x"83838383",
		1456 =>	x"85848383",
		1457 =>	x"83838383",
		1458 =>	x"83838383",
		1459 =>	x"83838383",
		1460 =>	x"85848383",
		1461 =>	x"83838383",
		1462 =>	x"83838383",
		1463 =>	x"83838383",
		1464 =>	x"85848383",
		1465 =>	x"83838383",
		1466 =>	x"83838383",
		1467 =>	x"83838E84",
		1468 =>	x"85848383",
		1469 =>	x"83838383",
		1470 =>	x"83838383",
		1471 =>	x"83838485",
		1472 =>	x"85848383", -- IMG_16x16_map_element_14
		1473 =>	x"83838383",
		1474 =>	x"83838383",
		1475 =>	x"83838485",
		1476 =>	x"848E8383",
		1477 =>	x"83838383",
		1478 =>	x"83838383",
		1479 =>	x"83838E84",
		1480 =>	x"83838383",
		1481 =>	x"83838383",
		1482 =>	x"83838383",
		1483 =>	x"83838383",
		1484 =>	x"83838383",
		1485 =>	x"83838383",
		1486 =>	x"83838383",
		1487 =>	x"83838383",
		1488 =>	x"83838383",
		1489 =>	x"83838383",
		1490 =>	x"83838383",
		1491 =>	x"83838383",
		1492 =>	x"83838383",
		1493 =>	x"83838383",
		1494 =>	x"83838383",
		1495 =>	x"83838383",
		1496 =>	x"83838383",
		1497 =>	x"83838383",
		1498 =>	x"83838383",
		1499 =>	x"83838383",
		1500 =>	x"83838383",
		1501 =>	x"83838383",
		1502 =>	x"83838383",
		1503 =>	x"83838383",
		1504 =>	x"83838383",
		1505 =>	x"83838383",
		1506 =>	x"83838383",
		1507 =>	x"83838383",
		1508 =>	x"83838383",
		1509 =>	x"83838383",
		1510 =>	x"83838383",
		1511 =>	x"83838383",
		1512 =>	x"83838383",
		1513 =>	x"83838383",
		1514 =>	x"83838383",
		1515 =>	x"83838383",
		1516 =>	x"83838383",
		1517 =>	x"83838383",
		1518 =>	x"83838383",
		1519 =>	x"83838383",
		1520 =>	x"83838383",
		1521 =>	x"83838383",
		1522 =>	x"83838383",
		1523 =>	x"83838383",
		1524 =>	x"83838383",
		1525 =>	x"83838383",
		1526 =>	x"83838383",
		1527 =>	x"83838383",
		1528 =>	x"84848484",
		1529 =>	x"84848484",
		1530 =>	x"84848484",
		1531 =>	x"84848484",
		1532 =>	x"85858585",
		1533 =>	x"85858585",
		1534 =>	x"85858585",
		1535 =>	x"85858585",
		1536 =>	x"85848383", -- IMG_16x16_map_element_15
		1537 =>	x"83838383",
		1538 =>	x"83838383",
		1539 =>	x"83838485",
		1540 =>	x"848E8383",
		1541 =>	x"83838383",
		1542 =>	x"83838383",
		1543 =>	x"83838485",
		1544 =>	x"83838383",
		1545 =>	x"83838383",
		1546 =>	x"83838383",
		1547 =>	x"83838485",
		1548 =>	x"83838383",
		1549 =>	x"83838383",
		1550 =>	x"83838383",
		1551 =>	x"83838485",
		1552 =>	x"83838383",
		1553 =>	x"83838383",
		1554 =>	x"83838383",
		1555 =>	x"83838485",
		1556 =>	x"83838383",
		1557 =>	x"83838383",
		1558 =>	x"83838383",
		1559 =>	x"83838485",
		1560 =>	x"83838383",
		1561 =>	x"83838383",
		1562 =>	x"83838383",
		1563 =>	x"83838485",
		1564 =>	x"83838383",
		1565 =>	x"83838383",
		1566 =>	x"83838383",
		1567 =>	x"83838485",
		1568 =>	x"83838383",
		1569 =>	x"83838383",
		1570 =>	x"83838383",
		1571 =>	x"83838485",
		1572 =>	x"83838383",
		1573 =>	x"83838383",
		1574 =>	x"83838383",
		1575 =>	x"83838485",
		1576 =>	x"83838383",
		1577 =>	x"83838383",
		1578 =>	x"83838383",
		1579 =>	x"83838485",
		1580 =>	x"83838383",
		1581 =>	x"83838383",
		1582 =>	x"83838383",
		1583 =>	x"83838485",
		1584 =>	x"83838383",
		1585 =>	x"83838383",
		1586 =>	x"83838383",
		1587 =>	x"83838485",
		1588 =>	x"83838383",
		1589 =>	x"83838383",
		1590 =>	x"83838383",
		1591 =>	x"83838485",
		1592 =>	x"848E8383",
		1593 =>	x"83838383",
		1594 =>	x"83838383",
		1595 =>	x"83838485",
		1596 =>	x"85848383",
		1597 =>	x"83838383",
		1598 =>	x"83838383",
		1599 =>	x"83838485",
		1600 =>	x"85848383", -- IMG_16x16_map_element_16
		1601 =>	x"83838383",
		1602 =>	x"83838383",
		1603 =>	x"83838485",
		1604 =>	x"85848383",
		1605 =>	x"83838383",
		1606 =>	x"83838383",
		1607 =>	x"83838485",
		1608 =>	x"85848383",
		1609 =>	x"83838383",
		1610 =>	x"83838383",
		1611 =>	x"83838485",
		1612 =>	x"85848383",
		1613 =>	x"83838383",
		1614 =>	x"83838383",
		1615 =>	x"83838485",
		1616 =>	x"85848383",
		1617 =>	x"83838383",
		1618 =>	x"83838383",
		1619 =>	x"83838485",
		1620 =>	x"85848383",
		1621 =>	x"83838383",
		1622 =>	x"83838383",
		1623 =>	x"83838485",
		1624 =>	x"85848383",
		1625 =>	x"83838383",
		1626 =>	x"83838383",
		1627 =>	x"83838485",
		1628 =>	x"85848383",
		1629 =>	x"83838383",
		1630 =>	x"83838383",
		1631 =>	x"83838485",
		1632 =>	x"85848383",
		1633 =>	x"83838383",
		1634 =>	x"83838383",
		1635 =>	x"83838485",
		1636 =>	x"85848383",
		1637 =>	x"83838383",
		1638 =>	x"83838383",
		1639 =>	x"83838485",
		1640 =>	x"85848383",
		1641 =>	x"83838383",
		1642 =>	x"83838383",
		1643 =>	x"83838485",
		1644 =>	x"85848383",
		1645 =>	x"83838383",
		1646 =>	x"83838383",
		1647 =>	x"83838485",
		1648 =>	x"85848383",
		1649 =>	x"83838383",
		1650 =>	x"83838383",
		1651 =>	x"83838485",
		1652 =>	x"85848383",
		1653 =>	x"83838383",
		1654 =>	x"83838383",
		1655 =>	x"83838485",
		1656 =>	x"85848383",
		1657 =>	x"83838383",
		1658 =>	x"83838383",
		1659 =>	x"83838485",
		1660 =>	x"85848383",
		1661 =>	x"83838383",
		1662 =>	x"83838383",
		1663 =>	x"83838485",
		1664 =>	x"85858585", -- IMG_16x16_map_element_17
		1665 =>	x"85858585",
		1666 =>	x"85858585",
		1667 =>	x"85858585",
		1668 =>	x"84848484",
		1669 =>	x"84848484",
		1670 =>	x"84848484",
		1671 =>	x"84848484",
		1672 =>	x"83838383",
		1673 =>	x"83838383",
		1674 =>	x"83838383",
		1675 =>	x"83838383",
		1676 =>	x"83838383",
		1677 =>	x"83838383",
		1678 =>	x"83838383",
		1679 =>	x"83838383",
		1680 =>	x"83838383",
		1681 =>	x"83838383",
		1682 =>	x"83838383",
		1683 =>	x"83838383",
		1684 =>	x"83838383",
		1685 =>	x"83838383",
		1686 =>	x"83838383",
		1687 =>	x"83838383",
		1688 =>	x"83838383",
		1689 =>	x"83838383",
		1690 =>	x"83838383",
		1691 =>	x"83838383",
		1692 =>	x"83838383",
		1693 =>	x"83838383",
		1694 =>	x"83838383",
		1695 =>	x"83838383",
		1696 =>	x"83838383",
		1697 =>	x"83838383",
		1698 =>	x"83838383",
		1699 =>	x"83838383",
		1700 =>	x"83838383",
		1701 =>	x"83838383",
		1702 =>	x"83838383",
		1703 =>	x"83838383",
		1704 =>	x"83838383",
		1705 =>	x"83838383",
		1706 =>	x"83838383",
		1707 =>	x"83838383",
		1708 =>	x"83838383",
		1709 =>	x"83838383",
		1710 =>	x"83838383",
		1711 =>	x"83838383",
		1712 =>	x"83838383",
		1713 =>	x"83838383",
		1714 =>	x"83838383",
		1715 =>	x"83838383",
		1716 =>	x"83838383",
		1717 =>	x"83838383",
		1718 =>	x"83838383",
		1719 =>	x"83838383",
		1720 =>	x"84848484",
		1721 =>	x"84848484",
		1722 =>	x"84848484",
		1723 =>	x"84848484",
		1724 =>	x"85858585",
		1725 =>	x"85858585",
		1726 =>	x"85858585",
		1727 =>	x"85858585",
		1728 =>	x"86878885", -- IMG_16x16_map_element_18
		1729 =>	x"85858585",
		1730 =>	x"85858585",
		1731 =>	x"85888786",
		1732 =>	x"898A8B8C",
		1733 =>	x"84848484",
		1734 =>	x"84848484",
		1735 =>	x"848F9087",
		1736 =>	x"888D8383",
		1737 =>	x"83838383",
		1738 =>	x"83838383",
		1739 =>	x"83838488",
		1740 =>	x"85848383",
		1741 =>	x"83838383",
		1742 =>	x"83838383",
		1743 =>	x"83838485",
		1744 =>	x"85848383",
		1745 =>	x"83838383",
		1746 =>	x"83838383",
		1747 =>	x"83838485",
		1748 =>	x"85848383",
		1749 =>	x"83838383",
		1750 =>	x"83838383",
		1751 =>	x"83838485",
		1752 =>	x"85848383",
		1753 =>	x"83838383",
		1754 =>	x"83838383",
		1755 =>	x"83838485",
		1756 =>	x"85848383",
		1757 =>	x"83838383",
		1758 =>	x"83838383",
		1759 =>	x"83838485",
		1760 =>	x"85848383",
		1761 =>	x"83838383",
		1762 =>	x"83838383",
		1763 =>	x"83838485",
		1764 =>	x"85848383",
		1765 =>	x"83838383",
		1766 =>	x"83838383",
		1767 =>	x"83838485",
		1768 =>	x"85848383",
		1769 =>	x"83838383",
		1770 =>	x"83838383",
		1771 =>	x"83838485",
		1772 =>	x"85848383",
		1773 =>	x"83838383",
		1774 =>	x"83838383",
		1775 =>	x"83838485",
		1776 =>	x"85848383",
		1777 =>	x"83838383",
		1778 =>	x"83838383",
		1779 =>	x"83838485",
		1780 =>	x"88848383",
		1781 =>	x"83838383",
		1782 =>	x"83838383",
		1783 =>	x"83838488",
		1784 =>	x"87908F84",
		1785 =>	x"84848484",
		1786 =>	x"84848484",
		1787 =>	x"848F9087",
		1788 =>	x"86878885",
		1789 =>	x"85858585",
		1790 =>	x"85858585",
		1791 =>	x"85888786",
		1792 =>	x"85858585", -- IMG_16x16_map_element_19
		1793 =>	x"85858585",
		1794 =>	x"85858585",
		1795 =>	x"85858585",
		1796 =>	x"84848484",
		1797 =>	x"84848484",
		1798 =>	x"84848484",
		1799 =>	x"84848484",
		1800 =>	x"83838383",
		1801 =>	x"83838383",
		1802 =>	x"83838383",
		1803 =>	x"83838383",
		1804 =>	x"83838383",
		1805 =>	x"83838383",
		1806 =>	x"83838383",
		1807 =>	x"83838383",
		1808 =>	x"83838383",
		1809 =>	x"83838383",
		1810 =>	x"83838383",
		1811 =>	x"83838383",
		1812 =>	x"83838383",
		1813 =>	x"83838383",
		1814 =>	x"83838383",
		1815 =>	x"83838383",
		1816 =>	x"83838383",
		1817 =>	x"83838383",
		1818 =>	x"83838383",
		1819 =>	x"83838383",
		1820 =>	x"83838383",
		1821 =>	x"83838383",
		1822 =>	x"83838383",
		1823 =>	x"83838383",
		1824 =>	x"83838383",
		1825 =>	x"83838383",
		1826 =>	x"83838383",
		1827 =>	x"83838383",
		1828 =>	x"83838383",
		1829 =>	x"83838383",
		1830 =>	x"83838383",
		1831 =>	x"83838383",
		1832 =>	x"83838383",
		1833 =>	x"83838383",
		1834 =>	x"83838383",
		1835 =>	x"83838383",
		1836 =>	x"83838383",
		1837 =>	x"83838383",
		1838 =>	x"83838383",
		1839 =>	x"83838383",
		1840 =>	x"83838383",
		1841 =>	x"83838383",
		1842 =>	x"83838383",
		1843 =>	x"83838383",
		1844 =>	x"83838383",
		1845 =>	x"83838383",
		1846 =>	x"83838383",
		1847 =>	x"83838383",
		1848 =>	x"83838383",
		1849 =>	x"83838383",
		1850 =>	x"83838383",
		1851 =>	x"83838383",
		1852 =>	x"83838383",
		1853 =>	x"83838383",
		1854 =>	x"83838383",
		1855 =>	x"83838383",
		1856 =>	x"85858585", -- IMG_16x16_map_element_20
		1857 =>	x"85858585",
		1858 =>	x"85858585",
		1859 =>	x"85888786",
		1860 =>	x"84848484",
		1861 =>	x"84848484",
		1862 =>	x"84848484",
		1863 =>	x"8C8B8A89",
		1864 =>	x"83838383",
		1865 =>	x"83838383",
		1866 =>	x"83838383",
		1867 =>	x"83838D88",
		1868 =>	x"83838383",
		1869 =>	x"83838383",
		1870 =>	x"83838383",
		1871 =>	x"83838485",
		1872 =>	x"83838383",
		1873 =>	x"83838383",
		1874 =>	x"83838383",
		1875 =>	x"83838485",
		1876 =>	x"83838383",
		1877 =>	x"83838383",
		1878 =>	x"83838383",
		1879 =>	x"83838485",
		1880 =>	x"83838383",
		1881 =>	x"83838383",
		1882 =>	x"83838383",
		1883 =>	x"83838485",
		1884 =>	x"83838383",
		1885 =>	x"83838383",
		1886 =>	x"83838383",
		1887 =>	x"83838485",
		1888 =>	x"83838383",
		1889 =>	x"83838383",
		1890 =>	x"83838383",
		1891 =>	x"83838485",
		1892 =>	x"83838383",
		1893 =>	x"83838383",
		1894 =>	x"83838383",
		1895 =>	x"83838485",
		1896 =>	x"83838383",
		1897 =>	x"83838383",
		1898 =>	x"83838383",
		1899 =>	x"83838485",
		1900 =>	x"83838383",
		1901 =>	x"83838383",
		1902 =>	x"83838383",
		1903 =>	x"83838485",
		1904 =>	x"83838383",
		1905 =>	x"83838383",
		1906 =>	x"83838383",
		1907 =>	x"83838485",
		1908 =>	x"83838383",
		1909 =>	x"83838383",
		1910 =>	x"83838383",
		1911 =>	x"83838485",
		1912 =>	x"83838383",
		1913 =>	x"83838383",
		1914 =>	x"83838383",
		1915 =>	x"83838485",
		1916 =>	x"83838383",
		1917 =>	x"83838383",
		1918 =>	x"83838383",
		1919 =>	x"83838485",
		1920 =>	x"86878885", -- IMG_16x16_map_element_21
		1921 =>	x"85858585",
		1922 =>	x"85858585",
		1923 =>	x"85858585",
		1924 =>	x"898A8B8C",
		1925 =>	x"84848484",
		1926 =>	x"84848484",
		1927 =>	x"84848484",
		1928 =>	x"888D8383",
		1929 =>	x"83838383",
		1930 =>	x"83838383",
		1931 =>	x"83838383",
		1932 =>	x"85848383",
		1933 =>	x"83838383",
		1934 =>	x"83838383",
		1935 =>	x"83838383",
		1936 =>	x"85848383",
		1937 =>	x"83838383",
		1938 =>	x"83838383",
		1939 =>	x"83838383",
		1940 =>	x"85848383",
		1941 =>	x"83838383",
		1942 =>	x"83838383",
		1943 =>	x"83838383",
		1944 =>	x"85848383",
		1945 =>	x"83838383",
		1946 =>	x"83838383",
		1947 =>	x"83838383",
		1948 =>	x"85848383",
		1949 =>	x"83838383",
		1950 =>	x"83838383",
		1951 =>	x"83838383",
		1952 =>	x"85848383",
		1953 =>	x"83838383",
		1954 =>	x"83838383",
		1955 =>	x"83838383",
		1956 =>	x"85848383",
		1957 =>	x"83838383",
		1958 =>	x"83838383",
		1959 =>	x"83838383",
		1960 =>	x"85848383",
		1961 =>	x"83838383",
		1962 =>	x"83838383",
		1963 =>	x"83838383",
		1964 =>	x"85848383",
		1965 =>	x"83838383",
		1966 =>	x"83838383",
		1967 =>	x"83838383",
		1968 =>	x"85848383",
		1969 =>	x"83838383",
		1970 =>	x"83838383",
		1971 =>	x"83838383",
		1972 =>	x"85848383",
		1973 =>	x"83838383",
		1974 =>	x"83838383",
		1975 =>	x"83838383",
		1976 =>	x"85848383",
		1977 =>	x"83838383",
		1978 =>	x"83838383",
		1979 =>	x"83838E84",
		1980 =>	x"85848383",
		1981 =>	x"83838383",
		1982 =>	x"83838383",
		1983 =>	x"83838485",
		1984 =>	x"86878885", -- IMG_16x16_map_element_22
		1985 =>	x"85858585",
		1986 =>	x"85858585",
		1987 =>	x"85888786",
		1988 =>	x"898A8B8C",
		1989 =>	x"84848484",
		1990 =>	x"84848484",
		1991 =>	x"8C8B8A89",
		1992 =>	x"888D8383",
		1993 =>	x"83838383",
		1994 =>	x"83838383",
		1995 =>	x"83838D88",
		1996 =>	x"85848383",
		1997 =>	x"83838383",
		1998 =>	x"83838383",
		1999 =>	x"83838485",
		2000 =>	x"85848383",
		2001 =>	x"83838383",
		2002 =>	x"83838383",
		2003 =>	x"83838485",
		2004 =>	x"85848383",
		2005 =>	x"83838383",
		2006 =>	x"83838383",
		2007 =>	x"83838485",
		2008 =>	x"85848383",
		2009 =>	x"83838383",
		2010 =>	x"83838383",
		2011 =>	x"83838485",
		2012 =>	x"85848383",
		2013 =>	x"83838383",
		2014 =>	x"83838383",
		2015 =>	x"83838485",
		2016 =>	x"85848383",
		2017 =>	x"83838383",
		2018 =>	x"83838383",
		2019 =>	x"83838485",
		2020 =>	x"85848383",
		2021 =>	x"83838383",
		2022 =>	x"83838383",
		2023 =>	x"83838485",
		2024 =>	x"85848383",
		2025 =>	x"83838383",
		2026 =>	x"83838383",
		2027 =>	x"83838485",
		2028 =>	x"85848383",
		2029 =>	x"83838383",
		2030 =>	x"83838383",
		2031 =>	x"83838485",
		2032 =>	x"85848383",
		2033 =>	x"83838383",
		2034 =>	x"83838383",
		2035 =>	x"83838485",
		2036 =>	x"85848383",
		2037 =>	x"83838383",
		2038 =>	x"83838383",
		2039 =>	x"83838485",
		2040 =>	x"85848383",
		2041 =>	x"83838383",
		2042 =>	x"83838383",
		2043 =>	x"83838485",
		2044 =>	x"85848383",
		2045 =>	x"83838383",
		2046 =>	x"83838383",
		2047 =>	x"83838485",
		2048 =>	x"85858585", -- IMG_16x16_map_element_23
		2049 =>	x"85858585",
		2050 =>	x"85858585",
		2051 =>	x"85888786",
		2052 =>	x"84848484",
		2053 =>	x"84848484",
		2054 =>	x"84848484",
		2055 =>	x"8C8B8A89",
		2056 =>	x"83838383",
		2057 =>	x"83838383",
		2058 =>	x"83838383",
		2059 =>	x"83838D88",
		2060 =>	x"83838383",
		2061 =>	x"83838383",
		2062 =>	x"83838383",
		2063 =>	x"83838485",
		2064 =>	x"83838383",
		2065 =>	x"83838383",
		2066 =>	x"83838383",
		2067 =>	x"83838485",
		2068 =>	x"83838383",
		2069 =>	x"83838383",
		2070 =>	x"83838383",
		2071 =>	x"83838485",
		2072 =>	x"83838383",
		2073 =>	x"83838383",
		2074 =>	x"83838383",
		2075 =>	x"83838485",
		2076 =>	x"83838383",
		2077 =>	x"83838383",
		2078 =>	x"83838383",
		2079 =>	x"83838485",
		2080 =>	x"83838383",
		2081 =>	x"83838383",
		2082 =>	x"83838383",
		2083 =>	x"83838485",
		2084 =>	x"83838383",
		2085 =>	x"83838383",
		2086 =>	x"83838383",
		2087 =>	x"83838485",
		2088 =>	x"83838383",
		2089 =>	x"83838383",
		2090 =>	x"83838383",
		2091 =>	x"83838485",
		2092 =>	x"83838383",
		2093 =>	x"83838383",
		2094 =>	x"83838383",
		2095 =>	x"83838485",
		2096 =>	x"83838383",
		2097 =>	x"83838383",
		2098 =>	x"83838383",
		2099 =>	x"83838485",
		2100 =>	x"83838383",
		2101 =>	x"83838383",
		2102 =>	x"83838383",
		2103 =>	x"83838485",
		2104 =>	x"848E8383",
		2105 =>	x"83838383",
		2106 =>	x"83838383",
		2107 =>	x"83838485",
		2108 =>	x"85848383",
		2109 =>	x"83838383",
		2110 =>	x"83838383",
		2111 =>	x"83838485",
		2112 =>	x"85848383", -- IMG_16x16_map_element_24
		2113 =>	x"83838383",
		2114 =>	x"83838383",
		2115 =>	x"83838383",
		2116 =>	x"85848383",
		2117 =>	x"83838383",
		2118 =>	x"83838383",
		2119 =>	x"83838383",
		2120 =>	x"85848383",
		2121 =>	x"83838383",
		2122 =>	x"83838383",
		2123 =>	x"83838383",
		2124 =>	x"85848383",
		2125 =>	x"83838383",
		2126 =>	x"83838383",
		2127 =>	x"83838383",
		2128 =>	x"85848383",
		2129 =>	x"83838383",
		2130 =>	x"83838383",
		2131 =>	x"83838383",
		2132 =>	x"85848383",
		2133 =>	x"83838383",
		2134 =>	x"83838383",
		2135 =>	x"83838383",
		2136 =>	x"85848383",
		2137 =>	x"83838383",
		2138 =>	x"83838383",
		2139 =>	x"83838383",
		2140 =>	x"85848383",
		2141 =>	x"83838383",
		2142 =>	x"83838383",
		2143 =>	x"83838383",
		2144 =>	x"85848383",
		2145 =>	x"83838383",
		2146 =>	x"83838383",
		2147 =>	x"83838383",
		2148 =>	x"85848383",
		2149 =>	x"83838383",
		2150 =>	x"83838383",
		2151 =>	x"83838383",
		2152 =>	x"85848383",
		2153 =>	x"83838383",
		2154 =>	x"83838383",
		2155 =>	x"83838383",
		2156 =>	x"85848383",
		2157 =>	x"83838383",
		2158 =>	x"83838383",
		2159 =>	x"83838383",
		2160 =>	x"85848383",
		2161 =>	x"83838383",
		2162 =>	x"83838383",
		2163 =>	x"83838383",
		2164 =>	x"85848383",
		2165 =>	x"83838383",
		2166 =>	x"83838383",
		2167 =>	x"83838383",
		2168 =>	x"85848383",
		2169 =>	x"83838383",
		2170 =>	x"83838383",
		2171 =>	x"83838383",
		2172 =>	x"85848383",
		2173 =>	x"83838383",
		2174 =>	x"83838383",
		2175 =>	x"83838383",
		2176 =>	x"83838383", -- IMG_16x16_map_element_25
		2177 =>	x"83838383",
		2178 =>	x"83838383",
		2179 =>	x"83838383",
		2180 =>	x"83838383",
		2181 =>	x"83838383",
		2182 =>	x"83838383",
		2183 =>	x"83838383",
		2184 =>	x"83838383",
		2185 =>	x"83838383",
		2186 =>	x"83838383",
		2187 =>	x"83838383",
		2188 =>	x"83838383",
		2189 =>	x"83838383",
		2190 =>	x"83838383",
		2191 =>	x"83838383",
		2192 =>	x"83838383",
		2193 =>	x"83838383",
		2194 =>	x"83838383",
		2195 =>	x"83838383",
		2196 =>	x"83838383",
		2197 =>	x"83838383",
		2198 =>	x"83838383",
		2199 =>	x"83838383",
		2200 =>	x"83838383",
		2201 =>	x"83838383",
		2202 =>	x"83838383",
		2203 =>	x"83838383",
		2204 =>	x"83838383",
		2205 =>	x"83838383",
		2206 =>	x"83838383",
		2207 =>	x"83838383",
		2208 =>	x"83838383",
		2209 =>	x"83838383",
		2210 =>	x"83838383",
		2211 =>	x"83838383",
		2212 =>	x"83838383",
		2213 =>	x"83838383",
		2214 =>	x"83838383",
		2215 =>	x"83838383",
		2216 =>	x"83838383",
		2217 =>	x"83838383",
		2218 =>	x"83838383",
		2219 =>	x"83838383",
		2220 =>	x"83838383",
		2221 =>	x"83838383",
		2222 =>	x"83838383",
		2223 =>	x"83838383",
		2224 =>	x"83838383",
		2225 =>	x"83838383",
		2226 =>	x"83838383",
		2227 =>	x"83838383",
		2228 =>	x"83838383",
		2229 =>	x"83838383",
		2230 =>	x"83838383",
		2231 =>	x"83838383",
		2232 =>	x"83838383",
		2233 =>	x"83838383",
		2234 =>	x"83838383",
		2235 =>	x"83838383",
		2236 =>	x"83838383",
		2237 =>	x"83838383",
		2238 =>	x"83838383",
		2239 =>	x"83838383",
		2240 =>	x"00000000", -- IMG_16x16_rock
		2241 =>	x"00000000",
		2242 =>	x"00000000",
		2243 =>	x"00000000",
		2244 =>	x"00000000",
		2245 =>	x"00000000",
		2246 =>	x"00000000",
		2247 =>	x"00000000",
		2248 =>	x"02030400",
		2249 =>	x"00000000",
		2250 =>	x"00000000",
		2251 =>	x"00000000",
		2252 =>	x"05060708",
		2253 =>	x"090A0506",
		2254 =>	x"07080B00",
		2255 =>	x"000C0D0E",
		2256 =>	x"0F101112",
		2257 =>	x"13141516",
		2258 =>	x"1718191A",
		2259 =>	x"1B1C1D0A",
		2260 =>	x"1E061F00",
		2261 =>	x"20062112",
		2262 =>	x"22232425",
		2263 =>	x"17102625",
		2264 =>	x"27062800",
		2265 =>	x"29062A00",
		2266 =>	x"2B062C00",
		2267 =>	x"2D062E00",
		2268 =>	x"2F063000",
		2269 =>	x"31063200",
		2270 =>	x"33063400",
		2271 =>	x"35063600",
		2272 =>	x"37063800",
		2273 =>	x"39063A00",
		2274 =>	x"07063B00",
		2275 =>	x"3C063D00",
		2276 =>	x"3E063F00",
		2277 =>	x"40064100",
		2278 =>	x"42064300",
		2279 =>	x"44064500",
		2280 =>	x"46064700",
		2281 =>	x"48064900",
		2282 =>	x"4A064B00",
		2283 =>	x"4C064D00",
		2284 =>	x"4E064F00",
		2285 =>	x"50065100",
		2286 =>	x"52065300",
		2287 =>	x"54065500",
		2288 =>	x"3C065600",
		2289 =>	x"57065800",
		2290 =>	x"57065900",
		2291 =>	x"57065A00",
		2292 =>	x"07080B00",
		2293 =>	x"5B5C5D5E",
		2294 =>	x"5F066000",
		2295 =>	x"61066200",
		2296 =>	x"63646566",
		2297 =>	x"6700680A",
		2298 =>	x"696A6B6C",
		2299 =>	x"6D0A0506",
		2300 =>	x"6E6F7071",
		2301 =>	x"72037323",
		2302 =>	x"74757616",
		2303 =>	x"77646378",
		2304 =>	x"79797979", -- IMG_16x16_smoke
		2305 =>	x"79797979",
		2306 =>	x"79797979",
		2307 =>	x"79797979",
		2308 =>	x"79797900",
		2309 =>	x"00000079",
		2310 =>	x"79797979",
		2311 =>	x"79000079",
		2312 =>	x"7979007B",
		2313 =>	x"7B7B0000",
		2314 =>	x"00000079",
		2315 =>	x"007B7B00",
		2316 =>	x"79007B7B",
		2317 =>	x"7B7B007B",
		2318 =>	x"7B7B7B79",
		2319 =>	x"007B7B00",
		2320 =>	x"7900007B",
		2321 =>	x"7B7B7B7B",
		2322 =>	x"7B7B7B00",
		2323 =>	x"7B7B7B00",
		2324 =>	x"7B7B7B7B",
		2325 =>	x"7B000000",
		2326 =>	x"7B7B0000",
		2327 =>	x"7B7B0079",
		2328 =>	x"7B7B7B7B",
		2329 =>	x"007B7B7B",
		2330 =>	x"007B7B7B",
		2331 =>	x"7B7B7B00",
		2332 =>	x"797B7B00",
		2333 =>	x"7B7B7B7B",
		2334 =>	x"0000007B",
		2335 =>	x"7B7B7B00",
		2336 =>	x"7B7B7B00",
		2337 =>	x"7B7B7B7B",
		2338 =>	x"7B7B007B",
		2339 =>	x"7B7B7B00",
		2340 =>	x"007B7B7B",
		2341 =>	x"7B7B7B7B",
		2342 =>	x"7B7B007B",
		2343 =>	x"7B7B7979",
		2344 =>	x"7B7B7B7B",
		2345 =>	x"7B7B7B7B",
		2346 =>	x"7B7B007B",
		2347 =>	x"00000079",
		2348 =>	x"79007B7B",
		2349 =>	x"7B7B7B7B",
		2350 =>	x"7B7B007B",
		2351 =>	x"7B7B7B79",
		2352 =>	x"79007B7B",
		2353 =>	x"7B7B7B7B",
		2354 =>	x"007B7B7B",
		2355 =>	x"7B7B0079",
		2356 =>	x"007B7B7B",
		2357 =>	x"7B007B7B",
		2358 =>	x"007B7B7B",
		2359 =>	x"7B7B0079",
		2360 =>	x"00000000",
		2361 =>	x"00007B7B",
		2362 =>	x"007B7B7B",
		2363 =>	x"7B000079",
		2364 =>	x"79797979",
		2365 =>	x"79790000",
		2366 =>	x"79790000",
		2367 =>	x"00797979",


--			***** MAP *****


		2368 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2369 =>	x"00000140", -- z: 0 rot: 0 ptr: 320
		2370 =>	x"00000180", -- z: 0 rot: 0 ptr: 384
		2371 =>	x"000001C0", -- z: 0 rot: 0 ptr: 448
		2372 =>	x"00000200", -- z: 0 rot: 0 ptr: 512
		2373 =>	x"00000240", -- z: 0 rot: 0 ptr: 576
		2374 =>	x"00000280", -- z: 0 rot: 0 ptr: 640
		2375 =>	x"000002C0", -- z: 0 rot: 0 ptr: 704
		2376 =>	x"00000300", -- z: 0 rot: 0 ptr: 768
		2377 =>	x"00000340", -- z: 0 rot: 0 ptr: 832
		2378 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2379 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2380 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2381 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2382 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2383 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2384 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2385 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2386 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2387 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2388 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2389 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2390 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2391 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2392 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2393 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2394 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2395 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2396 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2397 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2398 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2399 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2400 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2401 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2402 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2403 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2404 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2405 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2406 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2407 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2408 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2409 =>	x"00000380", -- z: 0 rot: 0 ptr: 896
		2410 =>	x"000003C0", -- z: 0 rot: 0 ptr: 960
		2411 =>	x"00000400", -- z: 0 rot: 0 ptr: 1024
		2412 =>	x"00000440", -- z: 0 rot: 0 ptr: 1088
		2413 =>	x"00000480", -- z: 0 rot: 0 ptr: 1152
		2414 =>	x"000004C0", -- z: 0 rot: 0 ptr: 1216
		2415 =>	x"00000500", -- z: 0 rot: 0 ptr: 1280
		2416 =>	x"00000540", -- z: 0 rot: 0 ptr: 1344
		2417 =>	x"00000580", -- z: 0 rot: 0 ptr: 1408
		2418 =>	x"000005C0", -- z: 0 rot: 0 ptr: 1472
		2419 =>	x"00000600", -- z: 0 rot: 0 ptr: 1536
		2420 =>	x"00000640", -- z: 0 rot: 0 ptr: 1600
		2421 =>	x"00000680", -- z: 0 rot: 0 ptr: 1664
		2422 =>	x"000006C0", -- z: 0 rot: 0 ptr: 1728
		2423 =>	x"00000700", -- z: 0 rot: 0 ptr: 1792
		2424 =>	x"00000740", -- z: 0 rot: 0 ptr: 1856
		2425 =>	x"000007C0", -- z: 0 rot: 0 ptr: 1984
		2426 =>	x"00000800", -- z: 0 rot: 0 ptr: 2048
		2427 =>	x"00000840", -- z: 0 rot: 0 ptr: 2112
		2428 =>	x"00000880", -- z: 0 rot: 0 ptr: 2176
		2429 =>	x"000004C0", -- z: 0 rot: 0 ptr: 1216
		2430 =>	x"00000600", -- z: 0 rot: 0 ptr: 1536
		2431 =>	x"000008C0", -- z: 0 rot: 0 ptr: 2240
		2432 =>	x"00000900", -- z: 0 rot: 0 ptr: 2304
		2433 =>	x"00000780", -- z: 0 rot: 0 ptr: 1920
		2434 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2435 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2436 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2437 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2438 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2439 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2440 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2441 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2442 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2443 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2444 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2445 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2446 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2447 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2448 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2449 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2450 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2451 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2452 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2453 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2454 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2455 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2456 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2457 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2458 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2459 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2460 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2461 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2462 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2463 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2464 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2465 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2466 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2467 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2468 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2469 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2470 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2471 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2472 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2473 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2474 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2475 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2476 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2477 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2478 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2479 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2480 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2481 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2482 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2483 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2484 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2485 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2486 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2487 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2488 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2489 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2490 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2491 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2492 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2493 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2494 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2495 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2496 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2497 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2498 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2499 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2500 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2501 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2502 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2503 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2504 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2505 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2506 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2507 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2508 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2509 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2510 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2511 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2512 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2513 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2514 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2515 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2516 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2517 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2518 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2519 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2520 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2521 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2522 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2523 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2524 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2525 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2526 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2527 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2528 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2529 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2530 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2531 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2532 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2533 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2534 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2535 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2536 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2537 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2538 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2539 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2540 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2541 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2542 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2543 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2544 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2545 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2546 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2547 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2548 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2549 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2550 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2551 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2552 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2553 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2554 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2555 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2556 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2557 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2558 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2559 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2560 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2561 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2562 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2563 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2564 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2565 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2566 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2567 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2568 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2569 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2570 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2571 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2572 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2573 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2574 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2575 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2576 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2577 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2578 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2579 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2580 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2581 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2582 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2583 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2584 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2585 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2586 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2587 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2588 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2589 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2590 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2591 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2592 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2593 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2594 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2595 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2596 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2597 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2598 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2599 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2600 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2601 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2602 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2603 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2604 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2605 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2606 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2607 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2608 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2609 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2610 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2611 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2612 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2613 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2614 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2615 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2616 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2617 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2618 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2619 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2620 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2621 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2622 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2623 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2624 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2625 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2626 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2627 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2628 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2629 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2630 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2631 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2632 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2633 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2634 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2635 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2636 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2637 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2638 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2639 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2640 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2641 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2642 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2643 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2644 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2645 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2646 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2647 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2648 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2649 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2650 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2651 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2652 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2653 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2654 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2655 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2656 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2657 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2658 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2659 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2660 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2661 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2662 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2663 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2664 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2665 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2666 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2667 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2668 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2669 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2670 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2671 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2672 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2673 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2674 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2675 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2676 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2677 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2678 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2679 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2680 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2681 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2682 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2683 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2684 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2685 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2686 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2687 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2688 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2689 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2690 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2691 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2692 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2693 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2694 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2695 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2696 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2697 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2698 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2699 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2700 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2701 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2702 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2703 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2704 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2705 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2706 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2707 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2708 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2709 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2710 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2711 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2712 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2713 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2714 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2715 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2716 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2717 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2718 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2719 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2720 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2721 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2722 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2723 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2724 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2725 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2726 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2727 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2728 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2729 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2730 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2731 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2732 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2733 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2734 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2735 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2736 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2737 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2738 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2739 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2740 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2741 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2742 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2743 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2744 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2745 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2746 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2747 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2748 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2749 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2750 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2751 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2752 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2753 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2754 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2755 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2756 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2757 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2758 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2759 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2760 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2761 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2762 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2763 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2764 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2765 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2766 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2767 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2768 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2769 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2770 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2771 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2772 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2773 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2774 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2775 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2776 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2777 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2778 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2779 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2780 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2781 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2782 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2783 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2784 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2785 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2786 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2787 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2788 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2789 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2790 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2791 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2792 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2793 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2794 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2795 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2796 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2797 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2798 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2799 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2800 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2801 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2802 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2803 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2804 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2805 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2806 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2807 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2808 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2809 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2810 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2811 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2812 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2813 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2814 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2815 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2816 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2817 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2818 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2819 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2820 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2821 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2822 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2823 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2824 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2825 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2826 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2827 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2828 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2829 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2830 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2831 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2832 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2833 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2834 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2835 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2836 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2837 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2838 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2839 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2840 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2841 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2842 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2843 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2844 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2845 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2846 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2847 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2848 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2849 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2850 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2851 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2852 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2853 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2854 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2855 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2856 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2857 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2858 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2859 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2860 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2861 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2862 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2863 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2864 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2865 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2866 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2867 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2868 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2869 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2870 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2871 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2872 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2873 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2874 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2875 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2876 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2877 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2878 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2879 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2880 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2881 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2882 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2883 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2884 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2885 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2886 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2887 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2888 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2889 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2890 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2891 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2892 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2893 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2894 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2895 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2896 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2897 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2898 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2899 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2900 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2901 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2902 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2903 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2904 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2905 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2906 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2907 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2908 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2909 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2910 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2911 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2912 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2913 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2914 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2915 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2916 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2917 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2918 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2919 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2920 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2921 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2922 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2923 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2924 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2925 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2926 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2927 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2928 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2929 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2930 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2931 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2932 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2933 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2934 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2935 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2936 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2937 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2938 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2939 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2940 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2941 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2942 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2943 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2944 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2945 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2946 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2947 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2948 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2949 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2950 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2951 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2952 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2953 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2954 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2955 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2956 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2957 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2958 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2959 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2960 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2961 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2962 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2963 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2964 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2965 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2966 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2967 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2968 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2969 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2970 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2971 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2972 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2973 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2974 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2975 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2976 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2977 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2978 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2979 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2980 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2981 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2982 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2983 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2984 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2985 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2986 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2987 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2988 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2989 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2990 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2991 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2992 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2993 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2994 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2995 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2996 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2997 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2998 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		2999 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3000 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3001 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3002 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3003 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3004 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3005 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3006 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3007 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3008 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3009 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3010 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3011 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3012 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3013 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3014 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3015 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3016 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3017 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3018 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3019 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3020 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3021 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3022 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3023 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3024 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3025 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3026 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3027 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3028 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3029 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3030 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3031 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3032 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3033 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3034 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3035 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3036 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3037 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3038 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3039 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3040 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3041 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3042 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3043 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3044 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3045 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3046 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3047 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3048 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3049 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3050 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3051 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3052 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3053 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3054 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3055 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3056 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3057 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3058 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3059 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3060 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3061 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3062 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3063 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3064 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3065 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3066 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3067 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3068 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3069 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3070 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3071 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3072 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3073 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3074 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3075 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3076 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3077 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3078 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3079 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3080 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3081 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3082 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3083 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3084 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3085 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3086 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3087 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3088 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3089 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3090 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3091 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3092 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3093 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3094 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3095 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3096 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3097 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3098 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3099 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3100 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3101 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3102 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3103 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3104 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3105 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3106 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3107 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3108 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3109 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3110 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3111 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3112 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3113 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3114 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3115 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3116 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3117 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3118 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3119 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3120 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3121 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3122 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3123 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3124 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3125 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3126 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3127 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3128 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3129 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3130 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3131 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3132 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3133 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3134 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3135 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3136 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3137 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3138 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3139 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3140 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3141 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3142 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3143 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3144 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3145 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3146 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3147 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3148 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3149 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3150 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3151 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3152 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3153 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3154 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3155 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3156 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3157 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3158 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3159 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3160 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3161 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3162 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3163 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3164 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3165 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3166 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3167 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3168 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3169 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3170 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3171 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3172 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3173 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3174 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3175 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3176 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3177 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3178 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3179 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3180 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3181 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3182 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3183 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3184 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3185 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3186 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3187 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3188 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3189 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3190 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3191 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3192 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3193 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3194 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3195 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3196 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3197 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3198 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3199 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3200 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3201 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3202 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3203 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3204 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3205 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3206 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3207 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3208 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3209 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3210 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3211 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3212 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3213 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3214 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3215 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3216 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3217 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3218 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3219 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3220 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3221 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3222 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3223 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3224 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3225 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3226 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3227 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3228 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3229 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3230 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3231 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3232 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3233 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3234 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3235 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3236 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3237 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3238 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3239 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3240 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3241 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3242 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3243 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3244 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3245 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3246 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3247 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3248 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3249 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3250 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3251 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3252 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3253 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3254 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3255 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3256 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3257 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3258 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3259 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3260 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3261 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3262 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3263 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3264 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3265 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3266 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3267 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3268 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3269 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3270 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3271 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3272 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3273 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3274 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3275 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3276 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3277 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3278 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3279 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3280 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3281 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3282 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3283 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3284 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3285 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3286 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3287 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3288 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3289 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3290 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3291 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3292 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3293 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3294 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3295 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3296 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3297 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3298 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3299 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3300 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3301 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3302 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3303 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3304 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3305 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3306 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3307 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3308 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3309 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3310 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3311 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3312 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3313 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3314 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3315 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3316 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3317 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3318 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3319 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3320 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3321 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3322 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3323 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3324 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3325 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3326 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3327 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3328 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3329 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3330 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3331 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3332 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3333 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3334 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3335 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3336 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3337 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3338 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3339 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3340 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3341 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3342 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3343 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3344 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3345 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3346 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3347 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3348 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3349 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3350 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3351 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3352 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3353 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3354 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3355 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3356 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3357 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3358 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3359 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3360 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3361 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3362 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3363 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3364 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3365 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3366 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3367 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3368 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3369 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3370 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3371 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3372 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3373 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3374 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3375 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3376 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3377 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3378 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3379 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3380 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3381 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3382 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3383 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3384 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3385 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3386 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3387 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3388 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3389 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3390 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3391 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3392 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3393 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3394 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3395 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3396 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3397 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3398 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3399 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3400 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3401 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3402 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3403 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3404 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3405 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3406 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3407 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3408 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3409 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3410 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3411 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3412 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3413 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3414 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3415 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3416 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3417 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3418 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3419 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3420 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3421 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3422 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3423 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3424 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3425 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3426 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3427 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3428 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3429 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3430 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3431 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3432 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3433 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3434 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3435 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3436 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3437 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3438 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3439 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3440 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3441 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3442 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3443 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3444 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3445 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3446 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3447 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3448 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3449 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3450 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3451 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3452 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3453 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3454 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3455 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3456 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3457 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3458 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3459 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3460 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3461 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3462 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3463 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3464 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3465 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3466 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3467 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3468 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3469 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3470 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3471 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3472 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3473 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3474 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3475 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3476 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3477 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3478 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3479 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3480 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3481 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3482 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3483 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3484 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3485 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3486 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3487 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3488 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3489 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3490 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3491 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3492 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3493 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3494 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3495 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3496 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3497 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3498 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3499 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3500 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3501 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3502 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3503 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3504 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3505 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3506 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3507 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3508 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3509 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3510 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3511 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3512 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3513 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3514 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3515 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3516 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3517 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3518 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3519 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3520 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3521 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3522 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3523 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3524 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3525 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3526 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3527 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3528 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3529 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3530 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3531 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3532 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3533 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3534 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3535 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3536 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3537 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3538 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3539 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3540 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3541 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3542 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3543 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3544 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3545 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3546 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3547 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3548 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3549 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3550 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3551 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3552 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3553 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3554 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3555 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3556 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3557 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3558 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3559 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3560 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3561 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3562 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3563 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3564 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3565 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3566 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3567 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3568 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3569 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3570 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3571 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3572 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3573 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3574 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3575 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3576 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3577 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3578 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3579 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3580 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3581 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3582 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3583 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3584 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3585 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3586 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3587 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3588 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3589 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3590 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3591 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3592 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3593 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3594 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3595 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3596 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3597 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3598 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3599 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3600 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3601 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3602 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3603 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3604 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3605 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3606 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3607 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3608 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3609 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3610 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3611 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3612 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3613 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3614 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3615 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3616 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3617 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3618 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3619 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3620 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3621 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3622 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3623 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3624 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3625 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3626 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3627 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3628 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3629 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3630 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3631 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3632 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3633 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3634 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3635 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3636 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3637 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		3638 =>	x"00000100", -- z: 0 rot: 0 ptr: 256
		others => x"00000000"
	);

begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;